module shifter_rotator(
	input logic[3:0] x,
	input logic[1:0] select,
	output logic[3:0] y
	);
//
endmodule