module mult_add(
	input logic [3:0] a0,
	input logic [3:0] a1,
	input logic [3:0] a2,
	input logic [3:0] a3,
	input logic [3:0] a4,
	input logic [3:0] a5,
	input logic [3:0] a6,
	input logic [3:0] a7,
	output logic [?:0] x);
//

endmodule