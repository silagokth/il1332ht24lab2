module mult_mnbit_tb #(parameter M = 4, parameter N = 4)(

);

//
endmodule